LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY FORWARD_UNIT IS
	PORT(
		Rs, Rt, EXMEM_Reg, MEMWB_Reg : IN STD_LOGIC_VECTOR(4 DOWNTO 0);
		EXMEM_RW, MEMWB_RW : IN STD_LOGIC; --REGISTER WRITE BACK CONTROL
		FWD_A, FWD_B : OUT STD_LOGIC_VECTOR(1 DOWNTO 0)
	);
END FORWARD_UNIT;

ARCHITECTURE Behaviour OF FORWARD_UNIT IS
BEGIN
	PROCESS(Rs, Rt)
	BEGIN
	No_Hazard:
		FWD_A <= "00";
		FWD_B <= "00";
	
	EX_Hazard:
		IF(EXMEM_RW = '1' AND
			EXMEM_Reg /= "00000" AND
			EXMEM_Reg = Rs)THEN
			FWD_A <= "10";
		END IF;
		
		IF(EXMEM_RW = '1' AND
			EXMEM_Reg /= "00000" AND
			EXMEM_Reg = Rt)THEN
			FWD_B <= "10";
		END IF;
		
	MEM_Hazard:
		IF(MEMWB_RW = '1' AND
			MEMWB_Reg /= "00000" AND
			NOT(EXMEM_RW = '1' AND EXMEM_Reg /= "00000" AND
			EXMEM_Reg = Rs) AND
			MEMWB_Reg = Rs) THEN
			FWD_A <= "01";
		END IF;
		
		IF(MEMWB_RW = '1' AND
			MEMWB_Reg /= "00000" AND
			NOT(EXMEM_RW = '1' AND EXMEM_Reg /= "00000" AND
			EXMEM_Reg = Rt) AND
			MEMWB_Reg = Rt) THEN
			FWD_B <= "01";
		END IF;
	END PROCESS;
END Behaviour;