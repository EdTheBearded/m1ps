LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY HAZARD_DETECTION IS
	PORT(
		IDEX_MemRead : IN STD_LOGIC;
		Rs, Rt, IDEX_Reg : IN STD_LOGIC_VECTOR(4 DOWNTO 0);
		PC_Wr, IFID_Wr, NOP : OUT STD_LOGIC
	);
END HAZARD_DETECTION;

ARCHITECTURE Behaviour OF HAZARD_DETECTION IS
BEGIN
	PROCESS(Rs, Rt)
	BEGIN
		IF(IDEX_MemRead = '1' AND
		  (IDEX_Reg = Rs OR IDEX_Reg = Rt)) THEN --Stall
			PC_Wr <= '0';
			IFID_Wr <= '0';
			NOP <= '0';
		ELSE --Don't Stall
			PC_Wr <= '1';
			IFID_Wr <= '1';
			NOP <= '1';
		END IF;
	END PROCESS;
END Behaviour;