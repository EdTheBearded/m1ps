LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY MUX4_1 IS
	PORT(
		IN0, IN1, IN2, IN3 : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		SEL : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
		CHOICE : OUT STD_LOGIC_VECTOR(31 DOWNTO 0)
	);
END MUX4_1;

ARCHITECTURE Behaviour OF MUX4_1 IS
BEGIN
	WITH SEL SELECT
		CHOICE <= IN0 WHEN "00",
				  IN1 WHEN "01",
				  IN2 WHEN "10",
				  IN3 WHEN OTHERS;
END Behaviour;