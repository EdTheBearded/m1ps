LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY MEMWB IS
	PORT(
		CLK, CLEAR : IN STD_LOGIC;
		ALUResult_I : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		INSTRUCTION_I : IN STD_LOGIC_VECTOR(4 DOWNTO 0);
		DMRead_I : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		MemToReg_I, Reg_Wr_I, Jal_In : IN STD_LOGIC;
		ALUResult_O : OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
		INSTRUCTION_O : OUT STD_LOGIC_VECTOR(4 DOWNTO 0);
		DMRead_O : OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
		MemToReg_O, Reg_Wr_O, Jal_Out : OUT STD_LOGIC
	);
END MEMWB;

ARCHITECTURE BEHAVIOUR OF MEMWB IS
BEGIN

	PROCESS(CLEAR, CLK)
	BEGIN
		IF CLEAR = '1' THEN
			ALUResult_O <= (OTHERS => '0');
			INSTRUCTION_O <= (OTHERS => '0');
			DMRead_O <= (OTHERS => '0');
			MemToReg_O <= '0';
			Reg_Wr_O <= '0';
			Jal_Out <= '0';
		ELSIF (CLK'EVENT AND CLK = '0') THEN
			ALUResult_O <= ALUResult_I;
			INSTRUCTION_O <= INSTRUCTION_I;
			DMRead_O <= DMRead_I;
			MemToReg_O <= MemToReg_I;
			Reg_Wr_O <= Reg_Wr_I;
			Jal_Out <= Jal_In;
		END IF;
	END PROCESS;
END BEHAVIOUR;