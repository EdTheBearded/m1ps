Library IEEE;
Use ieee.std_logic_1164.all;

ENTITY sign_ext IS
	PORT(
		immediate: IN STD_LOGIC_VECTOR(15 DOWNTO 0);
		ext_immediate: OUT STD_LOGIC_VECTOR(31 DOWNTO 0)
	);
END sign_ext;

ARCHITECTURE Behaviour OF sign_ext IS
BEGIN
	ext_immediate(31 DOWNTO 16) <= (OTHERS => immediate(15));
	ext_immediate(15 DOWNTO 0) <= immediate(15 DOWNTO 0);
END Behaviour;